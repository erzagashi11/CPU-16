`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.01.2024 02:28:53
// Design Name: 
// Module Name: MUX2IN1_16bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MUX2IN1_16bit(
    input [15:0] Hyrja0,
    input [15:0] Hyrja2,
    output [16:0] Dalja
    );
endmodule
